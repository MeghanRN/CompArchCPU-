`ifdef adder
`define adder

`endif //adder
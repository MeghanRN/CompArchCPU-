`ifdef clk
`define clk

`endif //clk
`include "mr_chips\components\alu.sv"
`include "mr_chips\components\clk.sv"
`include "mr_chips\components\decoder.sv"
`include "mr_chips\components\adder.sv"

`timescale 1ns/100ps


`ifdef decode
`define decode

`endif //decode
`include "mr_chips\mr_chips.sv"

`timescale 1ns/100ps


`include "mr_chips\components\alu.sv"
`include "mr_chips\components\clk.sv"
`include "mr_chips\components\decode.sv"
